library verilog;
use verilog.vl_types.all;
entity gaussian_blurrer_tf is
end gaussian_blurrer_tf;
