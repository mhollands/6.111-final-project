library verilog;
use verilog.vl_types.all;
entity main_fsm_tf is
end main_fsm_tf;
