library verilog;
use verilog.vl_types.all;
entity corner_detector_tf is
end corner_detector_tf;
