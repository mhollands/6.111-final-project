library verilog;
use verilog.vl_types.all;
entity sin_lookup_tf is
end sin_lookup_tf;
