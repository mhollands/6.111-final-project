library verilog;
use verilog.vl_types.all;
entity zbt_6111_sample is
    port(
        beep            : out    vl_logic;
        audio_reset_b   : out    vl_logic;
        ac97_sdata_out  : out    vl_logic;
        ac97_sdata_in   : in     vl_logic;
        ac97_synch      : out    vl_logic;
        ac97_bit_clock  : in     vl_logic;
        vga_out_red     : out    vl_logic_vector(7 downto 0);
        vga_out_green   : out    vl_logic_vector(7 downto 0);
        vga_out_blue    : out    vl_logic_vector(7 downto 0);
        vga_out_sync_b  : out    vl_logic;
        vga_out_blank_b : out    vl_logic;
        vga_out_pixel_clock: out    vl_logic;
        vga_out_hsync   : out    vl_logic;
        vga_out_vsync   : out    vl_logic;
        tv_out_ycrcb    : out    vl_logic_vector(9 downto 0);
        tv_out_reset_b  : out    vl_logic;
        tv_out_clock    : out    vl_logic;
        tv_out_i2c_clock: out    vl_logic;
        tv_out_i2c_data : out    vl_logic;
        tv_out_pal_ntsc : out    vl_logic;
        tv_out_hsync_b  : out    vl_logic;
        tv_out_vsync_b  : out    vl_logic;
        tv_out_blank_b  : out    vl_logic;
        tv_out_subcar_reset: out    vl_logic;
        tv_in_ycrcb     : in     vl_logic_vector(19 downto 0);
        tv_in_data_valid: in     vl_logic;
        tv_in_line_clock1: in     vl_logic;
        tv_in_line_clock2: in     vl_logic;
        tv_in_aef       : in     vl_logic;
        tv_in_hff       : in     vl_logic;
        tv_in_aff       : in     vl_logic;
        tv_in_i2c_clock : out    vl_logic;
        tv_in_i2c_data  : inout  vl_logic;
        tv_in_fifo_read : out    vl_logic;
        tv_in_fifo_clock: out    vl_logic;
        tv_in_iso       : out    vl_logic;
        tv_in_reset_b   : out    vl_logic;
        tv_in_clock     : out    vl_logic;
        ram0_data       : inout  vl_logic_vector(35 downto 0);
        ram0_address    : out    vl_logic_vector(18 downto 0);
        ram0_adv_ld     : out    vl_logic;
        ram0_clk        : out    vl_logic;
        ram0_cen_b      : out    vl_logic;
        ram0_ce_b       : out    vl_logic;
        ram0_oe_b       : out    vl_logic;
        ram0_we_b       : out    vl_logic;
        ram0_bwe_b      : out    vl_logic_vector(3 downto 0);
        ram1_data       : inout  vl_logic_vector(35 downto 0);
        ram1_address    : out    vl_logic_vector(18 downto 0);
        ram1_adv_ld     : out    vl_logic;
        ram1_clk        : out    vl_logic;
        ram1_cen_b      : out    vl_logic;
        ram1_ce_b       : out    vl_logic;
        ram1_oe_b       : out    vl_logic;
        ram1_we_b       : out    vl_logic;
        ram1_bwe_b      : out    vl_logic_vector(3 downto 0);
        clock_feedback_out: out    vl_logic;
        clock_feedback_in: in     vl_logic;
        flash_data      : inout  vl_logic_vector(15 downto 0);
        flash_address   : out    vl_logic_vector(23 downto 0);
        flash_ce_b      : out    vl_logic;
        flash_oe_b      : out    vl_logic;
        flash_we_b      : out    vl_logic;
        flash_reset_b   : out    vl_logic;
        flash_sts       : in     vl_logic;
        flash_byte_b    : out    vl_logic;
        rs232_txd       : out    vl_logic;
        rs232_rxd       : in     vl_logic;
        rs232_rts       : out    vl_logic;
        rs232_cts       : in     vl_logic;
        mouse_clock     : in     vl_logic;
        mouse_data      : in     vl_logic;
        keyboard_clock  : in     vl_logic;
        keyboard_data   : in     vl_logic;
        clock_27mhz     : in     vl_logic;
        clock1          : in     vl_logic;
        clock2          : in     vl_logic;
        disp_blank      : out    vl_logic;
        disp_data_out   : out    vl_logic;
        disp_clock      : out    vl_logic;
        disp_rs         : out    vl_logic;
        disp_ce_b       : out    vl_logic;
        disp_reset_b    : out    vl_logic;
        disp_data_in    : in     vl_logic;
        button0         : in     vl_logic;
        button1         : in     vl_logic;
        button2         : in     vl_logic;
        button3         : in     vl_logic;
        button_enter    : in     vl_logic;
        button_right    : in     vl_logic;
        button_left     : in     vl_logic;
        button_down     : in     vl_logic;
        button_up       : in     vl_logic;
        switch          : in     vl_logic_vector(7 downto 0);
        led             : out    vl_logic_vector(7 downto 0);
        user1           : inout  vl_logic_vector(31 downto 0);
        user2           : inout  vl_logic_vector(31 downto 0);
        user3           : inout  vl_logic_vector(31 downto 0);
        user4           : inout  vl_logic_vector(31 downto 0);
        daughtercard    : inout  vl_logic_vector(43 downto 0);
        systemace_data  : inout  vl_logic_vector(15 downto 0);
        systemace_address: out    vl_logic_vector(6 downto 0);
        systemace_ce_b  : out    vl_logic;
        systemace_we_b  : out    vl_logic;
        systemace_oe_b  : out    vl_logic;
        systemace_irq   : in     vl_logic;
        systemace_mpbrdy: in     vl_logic;
        analyzer1_data  : out    vl_logic_vector(15 downto 0);
        analyzer1_clock : out    vl_logic;
        analyzer2_data  : out    vl_logic_vector(15 downto 0);
        analyzer2_clock : out    vl_logic;
        analyzer3_data  : out    vl_logic_vector(15 downto 0);
        analyzer3_clock : out    vl_logic;
        analyzer4_data  : out    vl_logic_vector(15 downto 0);
        analyzer4_clock : out    vl_logic
    );
end zbt_6111_sample;
